.title KiCad schematic
.include "C:/AE/TLV1821/_models/BAT54.spice.txt"
.include "C:/AE/TLV1821/_models/tlv1821.lib"
R4 /VP /VOUT {RLOOP}
R5 /VP 0 {RREF}
XU1 /VP /VN VDD 0 /VOUT TLV1821
R6 VDD /VP {RPUP}
R3 VDD /VN {RPUN}
R2 /VDIV /VN {RIN2}
D1 0 /VDIV BAT54
V1 VDD 0 DC {VSUPPLY} 
V4 /VIN 0 DC SINE({Voffset} {Vamp} {Freq} {Td}) 
R1 /VIN /VDIV {RIN1}
.end
