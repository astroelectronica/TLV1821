.title KiCad schematic
.include "C:/AE/TLV1821/_models/c2012x7s2a105k125ae_p.mod"
.include "C:/AE/TLV1821/_models/tlv1821.lib"
R16 VCC /REF 100k
R14 VCC /COMMON {RDELAY}
XU4 /VIN /REF VCC 0 /COMMON TLV1821
XU5 /COMMON 0 C2012X7S2A105K125AE_p
V3 /VIN 0 PULSE({VL} {VH} {TD} {TR} {TF} {DUTY} {PERIODE} {NCYCLES})
R15 /REF 0 100k
XU3 /V3P /V3N VCC 0 /VOUT3 TLV1821
R12 VDD /VOUT3 100k
R11 /V3P /VOUT3 10Meg
R13 VCC /V3N 100k
XU2 /V2P /V2N VCC 0 /VOUT2 TLV1821
R5 /COMMON /V2P 10k
R9 /COMMON /V3P 10k
R7 /V2P /VOUT2 10Meg
R8 VDD /VOUT2 100k
R10 /V3N /V2N 51k
R1 /V1P /VOUT1 10Meg
R2 VDD /VOUT1 100k
R3 /V1N 0 51k
XU1 /V1P /V1N VCC 0 /VOUT1 TLV1821
R4 /COMMON /V1P 10k
R6 /V2N /V1N 51k
V2 VDD 0 DC {VLOGIC} 
V1 VCC 0 DC {VSUPPLY}
*
*qspice
*
*TLV1821
*Time delay generator
*AE01010821
*
*netlist
*.include TLV1821_delay.cir
*
*params
.param VSUPPLY=5
.param VLOGIC=3.3
.param RDELAY=100K
.param VL=0
.param VH=VSUPPLY
.param TD=10m
.param TR=50n
.param TF=50n
.param DUTY=150m
.param PERIODE=200m
.param NCYCLES=1
*
*transient response
.tran 0 200m 10n ;uic startup
* 
.end
